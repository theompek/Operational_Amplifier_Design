** Profile: "SCHEMATIC1-AcSweepAnalysisTemperature"  [ C:\ORCAD\Ergasia\ErgasiaTelestikou-PSpiceFiles\SCHEMATIC1\AcSweepAnalysisTemperature.sim ] 

** Creating circuit file "AcSweepAnalysisTemperature.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ergasiatelestikou-pspicefiles/nfet.lib" 
.LIB "../../../ergasiatelestikou-pspicefiles/pfet.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 400 0.1 1g
.TEMP 0 10 20 30 40 50 60 70
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
