** Profile: "SCHEMATIC1-SlewRateTemperature"  [ C:\ORCAD\Ergasia\ErgasiaTelestikou-PSpiceFiles\SCHEMATIC1\SlewRateTemperature.sim ] 

** Creating circuit file "SlewRateTemperature.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ergasiatelestikou-pspicefiles/nfet.lib" 
.LIB "../../../ergasiatelestikou-pspicefiles/pfet.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 3us 0 
.TEMP 0 10 20 30 40 50 60 70
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
